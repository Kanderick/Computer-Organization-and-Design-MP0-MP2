library verilog;
use verilog.vl_types.all;
entity add4 is
    generic(
        width           : integer := 32
    );
    port(
        a               : in     vl_logic_vector;
        f               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width : constant is 1;
end add4;
